library verilog;
use verilog.vl_types.all;
entity contador_assin_3_vlg_vec_tst is
end contador_assin_3_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity somadorcompleto_vlg_sample_tst is
    port(
        a1              : in     vl_logic;
        b1              : in     vl_logic;
        c               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end somadorcompleto_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity somadorcompleto_vlg_vec_tst is
end somadorcompleto_vlg_vec_tst;

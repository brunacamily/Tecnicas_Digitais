library verilog;
use verilog.vl_types.all;
entity exemplo8_vlg_vec_tst is
end exemplo8_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo12_vlg_vec_tst is
end exemplo12_vlg_vec_tst;

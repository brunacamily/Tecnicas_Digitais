library verilog;
use verilog.vl_types.all;
entity shifterESQ_vlg_vec_tst is
end shifterESQ_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity flip_flop_JK_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end flip_flop_JK_vlg_sample_tst;

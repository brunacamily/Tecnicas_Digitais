library verilog;
use verilog.vl_types.all;
entity exercicio2_vlg_check_tst is
    port(
        s               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end exercicio2_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity flip_flop_D_vlg_check_tst is
    port(
        saida           : in     vl_logic;
        saida_neg       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end flip_flop_D_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo1 is
    port(
        a               : in     vl_logic;
        b               : out    vl_logic
    );
end exemplo1;

library verilog;
use verilog.vl_types.all;
entity ff_jk_3bits_vlg_vec_tst is
end ff_jk_3bits_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo4_vlg_vec_tst is
end exemplo4_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo6_vlg_vec_tst is
end exemplo6_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo2_vlg_vec_tst is
end exemplo2_vlg_vec_tst;

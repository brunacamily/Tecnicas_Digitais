library verilog;
use verilog.vl_types.all;
entity exemplo3_vlg_vec_tst is
end exemplo3_vlg_vec_tst;

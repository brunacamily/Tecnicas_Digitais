library verilog;
use verilog.vl_types.all;
entity exercicio3_vlg_vec_tst is
end exercicio3_vlg_vec_tst;

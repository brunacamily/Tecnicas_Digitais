library verilog;
use verilog.vl_types.all;
entity xorSIMPLES_vlg_vec_tst is
end xorSIMPLES_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity somadorparalelo_vlg_vec_tst is
end somadorparalelo_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo5_vlg_vec_tst is
end exemplo5_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity bcd_ex3_vlg_vec_tst is
end bcd_ex3_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity xorSIMPLES_vlg_sample_tst is
    port(
        entrada01       : in     vl_logic;
        entrada02       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end xorSIMPLES_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity exercicio2_vlg_vec_tst is
end exercicio2_vlg_vec_tst;

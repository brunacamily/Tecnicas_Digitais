library verilog;
use verilog.vl_types.all;
entity somadorcompleto_vlg_check_tst is
    port(
        carry1          : in     vl_logic;
        sum1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end somadorcompleto_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo1_vlg_check_tst is
    port(
        b               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exemplo1_vlg_check_tst;

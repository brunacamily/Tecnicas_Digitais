library verilog;
use verilog.vl_types.all;
entity exemplo10_vlg_vec_tst is
end exemplo10_vlg_vec_tst;

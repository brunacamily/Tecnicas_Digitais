library verilog;
use verilog.vl_types.all;
entity muxPRINC_vlg_vec_tst is
end muxPRINC_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo7 is
    port(
        vetor           : in     vl_logic_vector(2 downto 0);
        s               : out    vl_logic
    );
end exemplo7;

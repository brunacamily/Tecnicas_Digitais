library verilog;
use verilog.vl_types.all;
entity exemplo15_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exemplo15_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity mux02_2x1_vlg_vec_tst is
end mux02_2x1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity xorSIMPLES_vlg_check_tst is
    port(
        Sout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end xorSIMPLES_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo7_vlg_vec_tst is
end exemplo7_vlg_vec_tst;

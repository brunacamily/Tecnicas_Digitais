library verilog;
use verilog.vl_types.all;
entity exercicio1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        ex3             : out    vl_logic_vector(3 downto 0)
    );
end exercicio1;

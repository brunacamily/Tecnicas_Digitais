library verilog;
use verilog.vl_types.all;
entity exercicio1_vlg_check_tst is
    port(
        ex3             : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end exercicio1_vlg_check_tst;

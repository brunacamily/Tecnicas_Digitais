library verilog;
use verilog.vl_types.all;
entity exemplo11_vlg_vec_tst is
end exemplo11_vlg_vec_tst;

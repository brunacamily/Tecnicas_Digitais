library verilog;
use verilog.vl_types.all;
entity reg_1bit_vlg_vec_tst is
end reg_1bit_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo1_vlg_vec_tst is
end exemplo1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo1_vlg_sample_tst is
    port(
        a               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end exemplo1_vlg_sample_tst;

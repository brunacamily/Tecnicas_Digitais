library verilog;
use verilog.vl_types.all;
entity cont_process_vlg_vec_tst is
end cont_process_vlg_vec_tst;

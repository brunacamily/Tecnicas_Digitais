library verilog;
use verilog.vl_types.all;
entity aula9_exemplo16_vlg_vec_tst is
end aula9_exemplo16_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo4_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exemplo4_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo9_vlg_vec_tst is
end exemplo9_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity exercicio1_vlg_vec_tst is
end exercicio1_vlg_vec_tst;

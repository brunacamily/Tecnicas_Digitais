library verilog;
use verilog.vl_types.all;
entity ff_jk_3bits_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ff_jk_3bits_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity exemplo15_vlg_vec_tst is
end exemplo15_vlg_vec_tst;

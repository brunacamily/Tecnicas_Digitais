library verilog;
use verilog.vl_types.all;
entity shifterDIR_vlg_vec_tst is
end shifterDIR_vlg_vec_tst;

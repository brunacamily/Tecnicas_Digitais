library verilog;
use verilog.vl_types.all;
entity Elogico_vlg_vec_tst is
end Elogico_vlg_vec_tst;

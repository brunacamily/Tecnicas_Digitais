library verilog;
use verilog.vl_types.all;
entity meiosomador_vlg_vec_tst is
end meiosomador_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity somadorparalelo2_vlg_vec_tst is
end somadorparalelo2_vlg_vec_tst;
